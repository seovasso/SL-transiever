`ifndef _const_vh_
`define _const_vh_

parameter APB_ADDR_WIDTH = 10;

//config reg width

//status reg width
parameter TX_STATUS_REG_WIDTH  = 1;
parameter RX_STATUS_REG_WIDTH  = 1;

//channel reg width


`endif
